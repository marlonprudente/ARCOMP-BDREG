library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bancoreg16bits is
	port(


	);
end entity;

architecture a_bancoreg16bits of bancoreg16bits is
	component reg16bits is
		port(

		);
	end component;